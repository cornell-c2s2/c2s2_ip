//================================================
// comb_float_divider.v
// 
// Combinational floating point multiplier
// Author: Mattie Lee (mll264)
// Additional credits: Barry Lyu (fl327), Xilai Dai (xd44)
//================================================

`ifndef COMB_FLOAT_DIVIDER_V
`define COMB_FLOAT_DIVIDER_V

module comb_float_divider #(
) (
  input  logic [31:0] in0,
  input  logic [31:0] in1,
  output logic [31:0] out
);

endmodule

`endif
