//SINE WAVE OF BIT_WIDTH = 32, DECIMAL_PT =  16
//FOR FFT OF SIZE = 128
`default_nettype none
module SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_128VRTL (
  output logic [32 - 1:0] sine_wave_out[0:128 - 1]
);
  assign sine_wave_out[0]   = 0;
  assign sine_wave_out[1]   = 3215;
  assign sine_wave_out[2]   = 6423;
  assign sine_wave_out[3]   = 9616;
  assign sine_wave_out[4]   = 12785;
  assign sine_wave_out[5]   = 15923;
  assign sine_wave_out[6]   = 19024;
  assign sine_wave_out[7]   = 22078;
  assign sine_wave_out[8]   = 25079;
  assign sine_wave_out[9]   = 28020;
  assign sine_wave_out[10]  = 30893;
  assign sine_wave_out[11]  = 33692;
  assign sine_wave_out[12]  = 36409;
  assign sine_wave_out[13]  = 39039;
  assign sine_wave_out[14]  = 41575;
  assign sine_wave_out[15]  = 44011;
  assign sine_wave_out[16]  = 46340;
  assign sine_wave_out[17]  = 48558;
  assign sine_wave_out[18]  = 50660;
  assign sine_wave_out[19]  = 52639;
  assign sine_wave_out[20]  = 54491;
  assign sine_wave_out[21]  = 56212;
  assign sine_wave_out[22]  = 57797;
  assign sine_wave_out[23]  = 59243;
  assign sine_wave_out[24]  = 60547;
  assign sine_wave_out[25]  = 61705;
  assign sine_wave_out[26]  = 62714;
  assign sine_wave_out[27]  = 63571;
  assign sine_wave_out[28]  = 64276;
  assign sine_wave_out[29]  = 64826;
  assign sine_wave_out[30]  = 65220;
  assign sine_wave_out[31]  = 65457;
  assign sine_wave_out[32]  = 65536;
  assign sine_wave_out[33]  = 65457;
  assign sine_wave_out[34]  = 65220;
  assign sine_wave_out[35]  = 64826;
  assign sine_wave_out[36]  = 64276;
  assign sine_wave_out[37]  = 63571;
  assign sine_wave_out[38]  = 62714;
  assign sine_wave_out[39]  = 61705;
  assign sine_wave_out[40]  = 60547;
  assign sine_wave_out[41]  = 59243;
  assign sine_wave_out[42]  = 57797;
  assign sine_wave_out[43]  = 56212;
  assign sine_wave_out[44]  = 54491;
  assign sine_wave_out[45]  = 52639;
  assign sine_wave_out[46]  = 50660;
  assign sine_wave_out[47]  = 48558;
  assign sine_wave_out[48]  = 46340;
  assign sine_wave_out[49]  = 44011;
  assign sine_wave_out[50]  = 41575;
  assign sine_wave_out[51]  = 39039;
  assign sine_wave_out[52]  = 36409;
  assign sine_wave_out[53]  = 33692;
  assign sine_wave_out[54]  = 30893;
  assign sine_wave_out[55]  = 28020;
  assign sine_wave_out[56]  = 25079;
  assign sine_wave_out[57]  = 22078;
  assign sine_wave_out[58]  = 19024;
  assign sine_wave_out[59]  = 15923;
  assign sine_wave_out[60]  = 12785;
  assign sine_wave_out[61]  = 9616;
  assign sine_wave_out[62]  = 6423;
  assign sine_wave_out[63]  = 3215;
  assign sine_wave_out[64]  = 0;
  assign sine_wave_out[65]  = -3215;
  assign sine_wave_out[66]  = -6423;
  assign sine_wave_out[67]  = -9616;
  assign sine_wave_out[68]  = -12785;
  assign sine_wave_out[69]  = -15923;
  assign sine_wave_out[70]  = -19024;
  assign sine_wave_out[71]  = -22078;
  assign sine_wave_out[72]  = -25079;
  assign sine_wave_out[73]  = -28020;
  assign sine_wave_out[74]  = -30893;
  assign sine_wave_out[75]  = -33692;
  assign sine_wave_out[76]  = -36409;
  assign sine_wave_out[77]  = -39039;
  assign sine_wave_out[78]  = -41575;
  assign sine_wave_out[79]  = -44011;
  assign sine_wave_out[80]  = -46340;
  assign sine_wave_out[81]  = -48558;
  assign sine_wave_out[82]  = -50660;
  assign sine_wave_out[83]  = -52639;
  assign sine_wave_out[84]  = -54491;
  assign sine_wave_out[85]  = -56212;
  assign sine_wave_out[86]  = -57797;
  assign sine_wave_out[87]  = -59243;
  assign sine_wave_out[88]  = -60547;
  assign sine_wave_out[89]  = -61705;
  assign sine_wave_out[90]  = -62714;
  assign sine_wave_out[91]  = -63571;
  assign sine_wave_out[92]  = -64276;
  assign sine_wave_out[93]  = -64826;
  assign sine_wave_out[94]  = -65220;
  assign sine_wave_out[95]  = -65457;
  assign sine_wave_out[96]  = -65536;
  assign sine_wave_out[97]  = -65457;
  assign sine_wave_out[98]  = -65220;
  assign sine_wave_out[99]  = -64826;
  assign sine_wave_out[100] = -64276;
  assign sine_wave_out[101] = -63571;
  assign sine_wave_out[102] = -62714;
  assign sine_wave_out[103] = -61705;
  assign sine_wave_out[104] = -60547;
  assign sine_wave_out[105] = -59243;
  assign sine_wave_out[106] = -57797;
  assign sine_wave_out[107] = -56212;
  assign sine_wave_out[108] = -54491;
  assign sine_wave_out[109] = -52639;
  assign sine_wave_out[110] = -50660;
  assign sine_wave_out[111] = -48558;
  assign sine_wave_out[112] = -46340;
  assign sine_wave_out[113] = -44011;
  assign sine_wave_out[114] = -41575;
  assign sine_wave_out[115] = -39039;
  assign sine_wave_out[116] = -36409;
  assign sine_wave_out[117] = -33692;
  assign sine_wave_out[118] = -30893;
  assign sine_wave_out[119] = -28020;
  assign sine_wave_out[120] = -25079;
  assign sine_wave_out[121] = -22078;
  assign sine_wave_out[122] = -19024;
  assign sine_wave_out[123] = -15923;
  assign sine_wave_out[124] = -12785;
  assign sine_wave_out[125] = -9616;
  assign sine_wave_out[126] = -6423;
  assign sine_wave_out[127] = -3215;
endmodule
