`ifndef SYSTOLICCTRL_V
`define SYSTOLICCTRL_V

module SystolicCtrl
#(
  parameter size = 16
)(
  input logic clk,
  input logic rst,
);



endmodule

`endif