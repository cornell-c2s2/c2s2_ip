// ===================================================================
// Author: Arjun Saini
// Date: 11/21/24
// Spec:  
// PARAMETERS --------------------------------------------------------
// 
// I/O ---------------------------------------------------------------
// - clk
// - reset
// ===================================================================

`ifndef LBIST_TOPLEVEL_V
`define LBIST_TOPLEVEL_V

module lbist_toplevel #(

  );

//============================LOCAL_PARAMETERS=================================

  
//================================DATAPATH=====================================


//===============================CTRL_LOGIC====================================


endmodule
`endif /* LBIST_TOPLEVEL_V */

