`ifndef fft_helpers_SINE_WAVE
`define fft_helpers_SINE_WAVE
`default_nettype none

// Macro to generate a sine table for N evenly spaced values from 0 to 2pi.
// Returns values in a fixedpoint format with D fractional bits and W total bits.
module fft_helpers_SineWave #(
  parameter int N = 8,
  parameter int W = 32,
  parameter int D = 16
) (
  output logic [W - 1:0] out[N]
);
  // Checks on parameters to make sure behavior is well defined.
  if (D >= 32) begin
    $error("D must be less than 32");
  end

  generate
    // arccos(-1) = pi
    real PI = $acos(-1);
    for (genvar i = 0; i < N; i++) begin
      real sinvalue = $sin(2 * PI * i / N);
      int  fixedptvalue = int'(sinvalue * 2.0 ** D);

      assign out[i] = {{(W - D - 1) {fixedptvalue[31]}}, fixedptvalue[D:0]};
    end
  endgenerate

endmodule

`endif
