//SINE WAVE OF BIT_WIDTH = 32, DECIMAL_PT =  16
//FOR FFT OF SIZE = 256
`default_nettype none
module SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_256VRTL (
  output logic [32 - 1:0] sine_wave_out[0:256 - 1]
);
  assign sine_wave_out[0]   = 0;
  assign sine_wave_out[1]   = 1608;
  assign sine_wave_out[2]   = 3215;
  assign sine_wave_out[3]   = 4821;
  assign sine_wave_out[4]   = 6423;
  assign sine_wave_out[5]   = 8022;
  assign sine_wave_out[6]   = 9616;
  assign sine_wave_out[7]   = 11204;
  assign sine_wave_out[8]   = 12785;
  assign sine_wave_out[9]   = 14359;
  assign sine_wave_out[10]  = 15923;
  assign sine_wave_out[11]  = 17479;
  assign sine_wave_out[12]  = 19024;
  assign sine_wave_out[13]  = 20557;
  assign sine_wave_out[14]  = 22078;
  assign sine_wave_out[15]  = 23586;
  assign sine_wave_out[16]  = 25079;
  assign sine_wave_out[17]  = 26557;
  assign sine_wave_out[18]  = 28020;
  assign sine_wave_out[19]  = 29465;
  assign sine_wave_out[20]  = 30893;
  assign sine_wave_out[21]  = 32302;
  assign sine_wave_out[22]  = 33692;
  assign sine_wave_out[23]  = 35061;
  assign sine_wave_out[24]  = 36409;
  assign sine_wave_out[25]  = 37736;
  assign sine_wave_out[26]  = 39039;
  assign sine_wave_out[27]  = 40319;
  assign sine_wave_out[28]  = 41575;
  assign sine_wave_out[29]  = 42806;
  assign sine_wave_out[30]  = 44011;
  assign sine_wave_out[31]  = 45189;
  assign sine_wave_out[32]  = 46340;
  assign sine_wave_out[33]  = 47464;
  assign sine_wave_out[34]  = 48558;
  assign sine_wave_out[35]  = 49624;
  assign sine_wave_out[36]  = 50660;
  assign sine_wave_out[37]  = 51665;
  assign sine_wave_out[38]  = 52639;
  assign sine_wave_out[39]  = 53581;
  assign sine_wave_out[40]  = 54491;
  assign sine_wave_out[41]  = 55368;
  assign sine_wave_out[42]  = 56212;
  assign sine_wave_out[43]  = 57022;
  assign sine_wave_out[44]  = 57797;
  assign sine_wave_out[45]  = 58538;
  assign sine_wave_out[46]  = 59243;
  assign sine_wave_out[47]  = 59913;
  assign sine_wave_out[48]  = 60547;
  assign sine_wave_out[49]  = 61144;
  assign sine_wave_out[50]  = 61705;
  assign sine_wave_out[51]  = 62228;
  assign sine_wave_out[52]  = 62714;
  assign sine_wave_out[53]  = 63162;
  assign sine_wave_out[54]  = 63571;
  assign sine_wave_out[55]  = 63943;
  assign sine_wave_out[56]  = 64276;
  assign sine_wave_out[57]  = 64571;
  assign sine_wave_out[58]  = 64826;
  assign sine_wave_out[59]  = 65043;
  assign sine_wave_out[60]  = 65220;
  assign sine_wave_out[61]  = 65358;
  assign sine_wave_out[62]  = 65457;
  assign sine_wave_out[63]  = 65516;
  assign sine_wave_out[64]  = 65536;
  assign sine_wave_out[65]  = 65516;
  assign sine_wave_out[66]  = 65457;
  assign sine_wave_out[67]  = 65358;
  assign sine_wave_out[68]  = 65220;
  assign sine_wave_out[69]  = 65043;
  assign sine_wave_out[70]  = 64826;
  assign sine_wave_out[71]  = 64571;
  assign sine_wave_out[72]  = 64276;
  assign sine_wave_out[73]  = 63943;
  assign sine_wave_out[74]  = 63571;
  assign sine_wave_out[75]  = 63162;
  assign sine_wave_out[76]  = 62714;
  assign sine_wave_out[77]  = 62228;
  assign sine_wave_out[78]  = 61705;
  assign sine_wave_out[79]  = 61144;
  assign sine_wave_out[80]  = 60547;
  assign sine_wave_out[81]  = 59913;
  assign sine_wave_out[82]  = 59243;
  assign sine_wave_out[83]  = 58538;
  assign sine_wave_out[84]  = 57797;
  assign sine_wave_out[85]  = 57022;
  assign sine_wave_out[86]  = 56212;
  assign sine_wave_out[87]  = 55368;
  assign sine_wave_out[88]  = 54491;
  assign sine_wave_out[89]  = 53581;
  assign sine_wave_out[90]  = 52639;
  assign sine_wave_out[91]  = 51665;
  assign sine_wave_out[92]  = 50660;
  assign sine_wave_out[93]  = 49624;
  assign sine_wave_out[94]  = 48558;
  assign sine_wave_out[95]  = 47464;
  assign sine_wave_out[96]  = 46340;
  assign sine_wave_out[97]  = 45189;
  assign sine_wave_out[98]  = 44011;
  assign sine_wave_out[99]  = 42806;
  assign sine_wave_out[100] = 41575;
  assign sine_wave_out[101] = 40319;
  assign sine_wave_out[102] = 39039;
  assign sine_wave_out[103] = 37736;
  assign sine_wave_out[104] = 36409;
  assign sine_wave_out[105] = 35061;
  assign sine_wave_out[106] = 33692;
  assign sine_wave_out[107] = 32302;
  assign sine_wave_out[108] = 30893;
  assign sine_wave_out[109] = 29465;
  assign sine_wave_out[110] = 28020;
  assign sine_wave_out[111] = 26557;
  assign sine_wave_out[112] = 25079;
  assign sine_wave_out[113] = 23586;
  assign sine_wave_out[114] = 22078;
  assign sine_wave_out[115] = 20557;
  assign sine_wave_out[116] = 19024;
  assign sine_wave_out[117] = 17479;
  assign sine_wave_out[118] = 15923;
  assign sine_wave_out[119] = 14359;
  assign sine_wave_out[120] = 12785;
  assign sine_wave_out[121] = 11204;
  assign sine_wave_out[122] = 9616;
  assign sine_wave_out[123] = 8022;
  assign sine_wave_out[124] = 6423;
  assign sine_wave_out[125] = 4821;
  assign sine_wave_out[126] = 3215;
  assign sine_wave_out[127] = 1608;
  assign sine_wave_out[128] = 0;
  assign sine_wave_out[129] = -1608;
  assign sine_wave_out[130] = -3215;
  assign sine_wave_out[131] = -4821;
  assign sine_wave_out[132] = -6423;
  assign sine_wave_out[133] = -8022;
  assign sine_wave_out[134] = -9616;
  assign sine_wave_out[135] = -11204;
  assign sine_wave_out[136] = -12785;
  assign sine_wave_out[137] = -14359;
  assign sine_wave_out[138] = -15923;
  assign sine_wave_out[139] = -17479;
  assign sine_wave_out[140] = -19024;
  assign sine_wave_out[141] = -20557;
  assign sine_wave_out[142] = -22078;
  assign sine_wave_out[143] = -23586;
  assign sine_wave_out[144] = -25079;
  assign sine_wave_out[145] = -26557;
  assign sine_wave_out[146] = -28020;
  assign sine_wave_out[147] = -29465;
  assign sine_wave_out[148] = -30893;
  assign sine_wave_out[149] = -32302;
  assign sine_wave_out[150] = -33692;
  assign sine_wave_out[151] = -35061;
  assign sine_wave_out[152] = -36409;
  assign sine_wave_out[153] = -37736;
  assign sine_wave_out[154] = -39039;
  assign sine_wave_out[155] = -40319;
  assign sine_wave_out[156] = -41575;
  assign sine_wave_out[157] = -42806;
  assign sine_wave_out[158] = -44011;
  assign sine_wave_out[159] = -45189;
  assign sine_wave_out[160] = -46340;
  assign sine_wave_out[161] = -47464;
  assign sine_wave_out[162] = -48558;
  assign sine_wave_out[163] = -49624;
  assign sine_wave_out[164] = -50660;
  assign sine_wave_out[165] = -51665;
  assign sine_wave_out[166] = -52639;
  assign sine_wave_out[167] = -53581;
  assign sine_wave_out[168] = -54491;
  assign sine_wave_out[169] = -55368;
  assign sine_wave_out[170] = -56212;
  assign sine_wave_out[171] = -57022;
  assign sine_wave_out[172] = -57797;
  assign sine_wave_out[173] = -58538;
  assign sine_wave_out[174] = -59243;
  assign sine_wave_out[175] = -59913;
  assign sine_wave_out[176] = -60547;
  assign sine_wave_out[177] = -61144;
  assign sine_wave_out[178] = -61705;
  assign sine_wave_out[179] = -62228;
  assign sine_wave_out[180] = -62714;
  assign sine_wave_out[181] = -63162;
  assign sine_wave_out[182] = -63571;
  assign sine_wave_out[183] = -63943;
  assign sine_wave_out[184] = -64276;
  assign sine_wave_out[185] = -64571;
  assign sine_wave_out[186] = -64826;
  assign sine_wave_out[187] = -65043;
  assign sine_wave_out[188] = -65220;
  assign sine_wave_out[189] = -65358;
  assign sine_wave_out[190] = -65457;
  assign sine_wave_out[191] = -65516;
  assign sine_wave_out[192] = -65536;
  assign sine_wave_out[193] = -65516;
  assign sine_wave_out[194] = -65457;
  assign sine_wave_out[195] = -65358;
  assign sine_wave_out[196] = -65220;
  assign sine_wave_out[197] = -65043;
  assign sine_wave_out[198] = -64826;
  assign sine_wave_out[199] = -64571;
  assign sine_wave_out[200] = -64276;
  assign sine_wave_out[201] = -63943;
  assign sine_wave_out[202] = -63571;
  assign sine_wave_out[203] = -63162;
  assign sine_wave_out[204] = -62714;
  assign sine_wave_out[205] = -62228;
  assign sine_wave_out[206] = -61705;
  assign sine_wave_out[207] = -61144;
  assign sine_wave_out[208] = -60547;
  assign sine_wave_out[209] = -59913;
  assign sine_wave_out[210] = -59243;
  assign sine_wave_out[211] = -58538;
  assign sine_wave_out[212] = -57797;
  assign sine_wave_out[213] = -57022;
  assign sine_wave_out[214] = -56212;
  assign sine_wave_out[215] = -55368;
  assign sine_wave_out[216] = -54491;
  assign sine_wave_out[217] = -53581;
  assign sine_wave_out[218] = -52639;
  assign sine_wave_out[219] = -51665;
  assign sine_wave_out[220] = -50660;
  assign sine_wave_out[221] = -49624;
  assign sine_wave_out[222] = -48558;
  assign sine_wave_out[223] = -47464;
  assign sine_wave_out[224] = -46340;
  assign sine_wave_out[225] = -45189;
  assign sine_wave_out[226] = -44011;
  assign sine_wave_out[227] = -42806;
  assign sine_wave_out[228] = -41575;
  assign sine_wave_out[229] = -40319;
  assign sine_wave_out[230] = -39039;
  assign sine_wave_out[231] = -37736;
  assign sine_wave_out[232] = -36409;
  assign sine_wave_out[233] = -35061;
  assign sine_wave_out[234] = -33692;
  assign sine_wave_out[235] = -32302;
  assign sine_wave_out[236] = -30893;
  assign sine_wave_out[237] = -29465;
  assign sine_wave_out[238] = -28020;
  assign sine_wave_out[239] = -26557;
  assign sine_wave_out[240] = -25079;
  assign sine_wave_out[241] = -23586;
  assign sine_wave_out[242] = -22078;
  assign sine_wave_out[243] = -20557;
  assign sine_wave_out[244] = -19024;
  assign sine_wave_out[245] = -17479;
  assign sine_wave_out[246] = -15923;
  assign sine_wave_out[247] = -14359;
  assign sine_wave_out[248] = -12785;
  assign sine_wave_out[249] = -11204;
  assign sine_wave_out[250] = -9616;
  assign sine_wave_out[251] = -8022;
  assign sine_wave_out[252] = -6423;
  assign sine_wave_out[253] = -4821;
  assign sine_wave_out[254] = -3215;
  assign sine_wave_out[255] = -1608;
endmodule
